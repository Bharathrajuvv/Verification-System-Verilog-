interface int_to(input bit clk,rst);
    logic  en;
  logic[3:0]  q;
endinterface
