interface int_to (input clk,rst);
  logic d;
  logic q;
endinterface

