interface add_if;
  logic  a,b,c;
  logic  sum,carry;
endinterface
