program test(add_if vif);
  environment env;
  initial begin
    env = new(vif);
    env.run();
  end
endprogram
