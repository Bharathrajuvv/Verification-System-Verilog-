Output:
Compiler version U-2023.03-SP2_Full64; Runtime version U-2023.03-SP2_Full64;  Aug 12 13:10 2025
__________ Driver _________
time=0 clk=0 rst=0 d=1 q=0
__________ Generator _________
time=10 clk=0 rst=0 d=1 q=0
__________ Monitor _________
time=10 clk=0 rst=0 d=1 q=0
__________ Driver _________
time=10 clk=0 rst=0 d=0 q=0
__________ Scoreboard _________
time=10 clk=0 rst=0 d=1 q=0
++++++++FAIL++++++++
__________ Generator _________
time=20 clk=0 rst=0 d=0 q=0
__________ Monitor _________
time=20 clk=0 rst=0 d=0 q=0
__________ Driver _________
time=20 clk=0 rst=0 d=1 q=0
__________ Scoreboard _________
time=20 clk=0 rst=0 d=0 q=0
++++++++PASS++++++++
__________ Generator _________
time=30 clk=0 rst=0 d=1 q=0
__________ Monitor _________
time=30 clk=0 rst=0 d=1 q=1
__________ Driver _________
time=30 clk=0 rst=0 d=1 q=0
__________ Scoreboard _________
time=30 clk=0 rst=0 d=1 q=1
++++++++PASS++++++++
__________ Generator _________
time=40 clk=0 rst=0 d=1 q=0
__________ Monitor _________
time=40 clk=0 rst=0 d=1 q=1
__________ Driver _________
time=40 clk=0 rst=0 d=0 q=0
__________ Scoreboard _________
time=40 clk=0 rst=0 d=1 q=1
++++++++PASS++++++++
__________ Generator _________
time=50 clk=0 rst=0 d=0 q=0
__________ Monitor _________
time=50 clk=0 rst=0 d=0 q=0
__________ Driver _________
time=50 clk=0 rst=0 d=0 q=0
__________ Scoreboard _________
time=50 clk=0 rst=0 d=0 q=0
++++++++PASS++++++++
__________ Generator _________
time=60 clk=0 rst=0 d=0 q=0
__________ Monitor _________
time=60 clk=0 rst=0 d=0 q=0
__________ Driver _________
time=60 clk=0 rst=0 d=1 q=0
__________ Scoreboard _________
time=60 clk=0 rst=0 d=0 q=0
++++++++PASS++++++++
__________ Generator _________
time=70 clk=0 rst=0 d=1 q=0
__________ Monitor _________
time=70 clk=0 rst=0 d=1 q=1
__________ Driver _________
time=70 clk=0 rst=0 d=1 q=0
__________ Scoreboard _________
time=70 clk=0 rst=0 d=1 q=1
++++++++PASS++++++++
__________ Generator _________
time=80 clk=0 rst=0 d=1 q=0
__________ Monitor _________
time=80 clk=0 rst=0 d=1 q=1
__________ Driver _________
time=80 clk=0 rst=0 d=0 q=0
__________ Scoreboard _________
time=80 clk=0 rst=0 d=1 q=1
++++++++PASS++++++++
__________ Generator _________
time=90 clk=0 rst=0 d=0 q=0
__________ Monitor _________
time=90 clk=0 rst=0 d=0 q=0
__________ Driver _________
time=90 clk=0 rst=0 d=0 q=0
__________ Scoreboard _________
time=90 clk=0 rst=0 d=0 q=0
++++++++PASS++++++++
__________ Generator _________
time=100 clk=0 rst=0 d=0 q=0
__________ Monitor _________
time=100 clk=0 rst=0 d=0 q=0
__________ Driver _________
time=100 clk=0 rst=0 d=0 q=0
__________ Scoreboard _________
time=100 clk=0 rst=0 d=0 q=0
++++++++PASS++++++++
__________ Generator _________
time=110 clk=0 rst=0 d=0 q=0
__________ Monitor _________
time=110 clk=0 rst=0 d=0 q=0
__________ Driver _________
time=110 clk=0 rst=0 d=0 q=0
__________ Scoreboard _________
time=110 clk=0 rst=0 d=0 q=0
++++++++PASS++++++++
__________ Generator _________
time=120 clk=0 rst=0 d=0 q=0
__________ Monitor _________
time=120 clk=0 rst=0 d=0 q=0
__________ Driver _________
time=120 clk=0 rst=0 d=1 q=0
__________ Scoreboard _________
time=120 clk=0 rst=0 d=0 q=0
++++++++PASS++++++++
__________ Generator _________
time=130 clk=0 rst=0 d=1 q=0
__________ Monitor _________
time=130 clk=0 rst=0 d=1 q=1
__________ Driver _________
time=130 clk=0 rst=0 d=0 q=0
__________ Scoreboard _________
time=130 clk=0 rst=0 d=1 q=1
++++++++PASS++++++++
__________ Generator _________
time=140 clk=0 rst=0 d=0 q=0
__________ Monitor _________
time=140 clk=0 rst=0 d=0 q=0
__________ Driver _________
time=140 clk=0 rst=0 d=0 q=0
__________ Scoreboard _________
time=140 clk=0 rst=0 d=0 q=0
++++++++PASS++++++++
__________ Generator _________
time=150 clk=0 rst=0 d=0 q=0
__________ Monitor _________
time=150 clk=0 rst=0 d=0 q=0
__________ Driver _________
time=150 clk=0 rst=0 d=0 q=0
__________ Scoreboard _________
time=150 clk=0 rst=0 d=0 q=0
++++++++PASS++++++++
__________ Generator _________
time=160 clk=0 rst=0 d=0 q=0
__________ Monitor _________
time=160 clk=0 rst=0 d=0 q=0
__________ Scoreboard _________
time=160 clk=0 rst=0 d=0 q=0
++++++++PASS++++++++
$finish called from file "testbench.sv", line 17.
$finish at simulation time                  210

